--------------------------------------------------------%
-- ULA                                                  %
-- Entradas: a, b e c                                   %
-- Saidas: saida, soma e carry                          %
-- Dependencias: meiosomador.vhd                        %
--------------------------------------------------------% 